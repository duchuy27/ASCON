module tb_spi_top();
    parameter MAIN_CLK_DELAY = 2;  // 25 MHz

    logic r_Rst_L     = 1'b0;  
    logic w_SPI_Clk;
    logic r_Clk       = 1'b0;
    logic w_SPI_MOSI;

    // Master Specific
    logic [7:0] r_Master_TX_Byte = 0;
    logic r_Master_TX_DV = 1'b0;
    logic w_Master_TX_Ready;
    logic r_Master_RX_DV;
    logic [7:0] r_Master_RX_Byte;

    // Clock Generators:
    always #(MAIN_CLK_DELAY) r_Clk = ~r_Clk;

    // Instantiate the spi_top module
    spi_top dut (
        // Control/Data Signals,
        .i_Rst_L(r_Rst_L),     // FPGA Reset
        .i_Clk(r_Clk),         // FPGA Clock
        
        // TX (MOSI) Signals
        .i_TX_Byte(r_Master_TX_Byte),     // Byte to transmit on MOSI
        .i_TX_DV(r_Master_TX_DV),         // Data Valid Pulse with i_TX_Byte
        .o_TX_Ready(w_Master_TX_Ready),   // Transmit Ready for Byte
        
        // RX (MISO) Signals
        .o_RX_DV(r_Master_RX_DV),       // Data Valid pulse (1 clock cycle)
        .o_RX_Byte(r_Master_RX_Byte),   // Byte received on MISO

        // SPI Interface
        .o_SPI_Clk(w_SPI_Clk),
        .i_SPI_MISO(w_SPI_MOSI),
        .o_SPI_MOSI(w_SPI_MOSI)
    );

    // Reset generation
    initial begin
        r_Rst_L = 0;
        #10;
        r_Rst_L = 1;
    end

    // Test sequence
    initial begin
        // Required for EDA Playground
        $dumpfile("dump.vcd"); 
        $dumpvars;

        // Wait for reset to settle
        #20;

        // Test single byte
        r_Master_TX_DV = 1'b1;
        r_Master_TX_Byte = 8'hC1;
        #10;

        if (w_Master_TX_Ready) begin
            r_Master_TX_Byte = 8'hA2;
            #10;
        end
        
        if (w_Master_TX_Ready) begin
            r_Master_TX_Byte = 8'hB3;
            #10;
        end
        $display("Sent out 0xC1, Received 0x%X", r_Master_RX_Byte);

        // Finish simulation
        #10;
        $finish();
    end
endmodule
